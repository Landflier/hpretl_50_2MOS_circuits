** sch_path: /home/vasil/CAD_VLSI/analog-circuit-design/xschem/dc_lv_nmos.sch
**.subckt dc_lv_nmos
Vgs net1 GND 0.65
Vds net3 GND 1.5
XM1 net2 net1 GND GND sg13_lv_nmos w=1.3u l=0.13u ng=1 m=1
Vd net3 net2 0
.save i(vd)
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.temp 27
.control
save all
save @n.xm1.nsg13_lv_nmos[gm]
save @n.xm1.nsg13_lv_nmos[gds]
save @n.xm1.nsg13_lv_nmos[vth]
save @n.xm1.nsg13_lv_nmos[cgg]
save @n.xm1.nsg13_lv_nmos[cgd]
save @n.xm1.nsg13_lv_nmos[vdss]
save @n.xm1.nsg13_lv_nmos[fug]
save @n.xm1.nsg13_lv_nmos[rg]
save @n.xm1.nsg13_lv_nmos[sid]
op
write dc_lv_nmos.raw
set appendwrite
dc Vds 0 1.5 0.01 Vgs 0 1.5 0.1
write dc_lv_nmos.raw
quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
